module And (
    input a, b;
    output out
);
  nand n1(a, b, out);

endmodule